module reg65(outputs, in, clk);
    input [64:0] in;
    input clk;
    output [64:0] outputs;
    wire in_en, reset;
    assign in_en = 1'b1;
    assign reset = 1'b0;

    dffe_ref reg0(outputs[0], in[0], clk, in_en, reset);
    dffe_ref reg1(outputs[1], in[1], clk, in_en, reset);
    dffe_ref reg2(outputs[2], in[2], clk, in_en, reset);
    dffe_ref reg3(outputs[3], in[3], clk, in_en, reset);
    dffe_ref reg4(outputs[4], in[4], clk, in_en, reset);
    dffe_ref reg5(outputs[5], in[5], clk, in_en, reset);
    dffe_ref reg6(outputs[6], in[6], clk, in_en, reset);
    dffe_ref reg7(outputs[7], in[7], clk, in_en, reset);
    dffe_ref reg8(outputs[8], in[8], clk, in_en, reset);
    dffe_ref reg9(outputs[9], in[9], clk, in_en, reset);
    dffe_ref reg10(outputs[10], in[10], clk, in_en, reset);
    dffe_ref reg11(outputs[11], in[11], clk, in_en, reset);
    dffe_ref reg12(outputs[12], in[12], clk, in_en, reset);
    dffe_ref reg13(outputs[13], in[13], clk, in_en, reset);
    dffe_ref reg14(outputs[14], in[14], clk, in_en, reset);
    dffe_ref reg15(outputs[15], in[15], clk, in_en, reset);
    dffe_ref reg16(outputs[16], in[16], clk, in_en, reset);
    dffe_ref reg17(outputs[17], in[17], clk, in_en, reset);
    dffe_ref reg18(outputs[18], in[18], clk, in_en, reset);
    dffe_ref reg19(outputs[19], in[19], clk, in_en, reset);
    dffe_ref reg20(outputs[20], in[20], clk, in_en, reset);
    dffe_ref reg21(outputs[21], in[21], clk, in_en, reset);
    dffe_ref reg22(outputs[22], in[22], clk, in_en, reset);
    dffe_ref reg23(outputs[23], in[23], clk, in_en, reset);
    dffe_ref reg24(outputs[24], in[24], clk, in_en, reset);
    dffe_ref reg25(outputs[25], in[25], clk, in_en, reset);
    dffe_ref reg26(outputs[26], in[26], clk, in_en, reset);
    dffe_ref reg27(outputs[27], in[27], clk, in_en, reset);
    dffe_ref reg28(outputs[28], in[28], clk, in_en, reset);
    dffe_ref reg29(outputs[29], in[29], clk, in_en, reset);
    dffe_ref reg30(outputs[30], in[30], clk, in_en, reset);
    dffe_ref reg31(outputs[31], in[31], clk, in_en, reset);
    dffe_ref reg32(outputs[32], in[32], clk, in_en, reset);
    dffe_ref reg33(outputs[33], in[33], clk, in_en, reset);
    dffe_ref reg34(outputs[34], in[34], clk, in_en, reset);
    dffe_ref reg35(outputs[35], in[35], clk, in_en, reset);
    dffe_ref reg36(outputs[36], in[36], clk, in_en, reset);
    dffe_ref reg37(outputs[37], in[37], clk, in_en, reset);
    dffe_ref reg38(outputs[38], in[38], clk, in_en, reset);
    dffe_ref reg39(outputs[39], in[39], clk, in_en, reset);
    dffe_ref reg40(outputs[40], in[40], clk, in_en, reset);
    dffe_ref reg41(outputs[41], in[41], clk, in_en, reset);
    dffe_ref reg42(outputs[42], in[42], clk, in_en, reset);
    dffe_ref reg43(outputs[43], in[43], clk, in_en, reset);
    dffe_ref reg44(outputs[44], in[44], clk, in_en, reset);
    dffe_ref reg45(outputs[45], in[45], clk, in_en, reset);
    dffe_ref reg46(outputs[46], in[46], clk, in_en, reset);
    dffe_ref reg47(outputs[47], in[47], clk, in_en, reset);
    dffe_ref reg48(outputs[48], in[48], clk, in_en, reset);
    dffe_ref reg49(outputs[49], in[49], clk, in_en, reset);
    dffe_ref reg50(outputs[50], in[50], clk, in_en, reset);
    dffe_ref reg51(outputs[51], in[51], clk, in_en, reset);
    dffe_ref reg52(outputs[52], in[52], clk, in_en, reset);
    dffe_ref reg53(outputs[53], in[53], clk, in_en, reset);
    dffe_ref reg54(outputs[54], in[54], clk, in_en, reset);
    dffe_ref reg55(outputs[55], in[55], clk, in_en, reset);
    dffe_ref reg56(outputs[56], in[56], clk, in_en, reset);
    dffe_ref reg57(outputs[57], in[57], clk, in_en, reset);
    dffe_ref reg58(outputs[58], in[58], clk, in_en, reset);
    dffe_ref reg59(outputs[59], in[59], clk, in_en, reset);
    dffe_ref reg60(outputs[60], in[60], clk, in_en, reset);
    dffe_ref reg61(outputs[61], in[61], clk, in_en, reset);
    dffe_ref reg62(outputs[62], in[62], clk, in_en, reset);
    dffe_ref reg63(outputs[63], in[63], clk, in_en, reset);
    dffe_ref reg64(outputs[64], in[64], clk, in_en, reset);

endmodule